module ALUControl(
    output [3:0] mode,
    input op,
    input [5:0] func
);
    assign mode = 0;
endmodule