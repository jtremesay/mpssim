module Control(
    output dr_sel, jump, branch, mem_to_reg, alu_op, mem_write, alu_sel, dr_write,
    input [5:0] op
);

endmodule