module Adder(output [31:0] z, input [31:0] a, b);
    assign z = a + b;
endmodule